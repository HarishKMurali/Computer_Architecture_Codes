`include "fp_multiplier.v"

module top;

	reg [31:0]a, b;
	reg clk;
	wire [31:0]out;
	initial begin
		clk=0;
	end

	always 
		#1 clk=~clk;

	fp_multiplier FP1 (a, b, out,clk);

	initial
	begin

		//+ve,+ve
		 a=32'b0_10001000_11101100000101000000100;	// 984.156494140625
		 b=32'b0_10001011_01101110110100100101010;	// 5869.1455078125

		 //#30 a = 32'b0_10000000_11110000000000000000000;b = 32'b1_10000000_11000000000000000000000;		// 3.5

		//#5 $display("A:\t %b %b %b\nB:\t %b %b %b\noutput:\t %b %b %b\n", a[31], a[30:23], a[22:0], b[31], b[30:23], b[22:0], out[31], out[30:23], out[22:0]);
		//==> 32'b0 10010101 01100000100011000111011
		#35 $finish();
	// 	//+ve,-ve
	// 	#10 a = 32'b0_10000000_11110000000000000000000;		// 3.875
	// 	#10 b = 32'b1_10000000_11000000000000000000000;		// 3.5
	// 	#10 $display("A:\t %b %b %b\nB:\t %b %b %b\noutput:\t %b %b %b\n", a[31], a[30:23], a[22:0], b[31], b[30:23], b[22:0], out[31], out[30:23], out[22:0]);
	// // ==> 32'b1 10000010 10110010000000000000000 

	// 	#5 a=32'b1_10001011_00000100010111100100111;	// -4165.89404296875
	// 	#5 b=32'b0_10000110_00111000011000001110111;	// 156.18931579589844
	// 	#5 $display("A:\t %b %b %b\nB:\t %b %b %b\noutput:\t %b %b %b\n", a[31], a[30:23], a[22:0], b[31], b[30:23], b[22:0], out[31], out[30:23], out[22:0]);
		
	// 	//zero*number
	// 	#15 a = 32'b0_00000000_00000000000000000000000;		// 3.875
	// 	#15 b = 32'b0_10000000_00000000000000000000000;		// 3.5
	// 	#15 $display("A:\t %b %b %b\nB:\t %b %b %b\noutput:\t %b %b %b\n", a[31], a[30:23], a[22:0], b[31], b[30:23], b[22:0], out[31], out[30:23], out[22:0]);

	// 	//zero * inf
	// 	#20 a = 32'b0_00000000_00000000000000000000000;		// zero
	// 	#20 b = 32'b0_11111111_00000000000000000000000;		// infinity
	// 	#20 $display("A:\t %b %b %b\nB:\t %b %b %b\noutput:\t %b %b %b\n", a[31], a[30:23], a[22:0], b[31], b[30:23], b[22:0], out[31], out[30:23], out[22:0]);
		
	// 	//inf * inf
	// 	#20 a = 32'b0_11111111_00000000000000000000000;		// zero
	// 	#20 b = 32'b0_11111111_00000000000000000000000;		// infinity
	// 	#20 $display("A:\t %b %b %b\nB:\t %b %b %b\noutput:\t %b %b %b\n", a[31], a[30:23], a[22:0], b[31], b[30:23], b[22:0], out[31], out[30:23], out[22:0]);
	// 	// a=32'b1_10001100_10010101011110010100000;	// -12975.15625
	// 	// b=32'b1_10001110_01101111000011000110000;	// -46982.1875
		// #5 $display("%b_%b_%b", out[31], out[30:23], out[22:0]);

	end
	initial 
        $monitor($time,"A = %b, B = %b,out= %b",a,b,out);

endmodule