`include "FP_adder.v"

module FP_adder_tb;
reg [31:0]a, b;
wire [31:0]out;

FP_adder FP1 (a, b, out);

initial
begin

	//a=32'b0_10001011_11110100000000000000000; //8000
	//b=32'b1_10001011_01110111000000000000000; //-6000
	// +ve +ve 
	//a = 32'b0_10000000_11110000000000000000000;		// 3.875
	//b = 32'b0_10000000_11000000000000000000000;		// 3.5
	// ==> 32'b0_10000001_11011000000000000000000  ans = 7.375

	//-ve +ve
	//a = 32'b1_10000000_11100000000000000000000;		// -3.75
	//b = 32'b0_10000000_11000000000000000000000;		// 3.5 // ans:1 01111101 00000000000000000000000
	
	// -ve -ve
	// a =	32'b1_10000010_00111000000000000000000;
	// b =	32'b1_10000010_00111000000000000000000;

	// a = 32'b0_10000010_00111000000000000000000;
	// b = 32'b0_10000000_11000000000000000000000;
	
	// infinity case(+,-)
	// a = 32'b0_11111111_00000000000000000000000;
	// b = 32'b1_11111100_00000000000000000000000;

	// infinity case(+,+)
	a = 32'b0_11111111_00000000000000000000000;
	 b = 32'b0_11111111_00000000000000000000000;

	//+ve -ve
	// a = 32'b0_01111110_01100000000000000000000;
	// b = 32'b1_01111110_00100000000000000000000;// ans:0 01111100 00000000000000000000000

	// b = 32'b0_01111111_00000000000000000000000;
	 //a = 32'h0000;
	//b = 32'h0000;
	#5 $display("A:\t %b %b %b", a[31], a[30:23], a[22:0]);
	#5 $display("B:\t %b %b %b", b[31], b[30:23], b[22:0]);
	#5 $display("output:\t %b %b %b", out[31], out[30:23], out[22:0]);
end


endmodule