module mux(a,b,s,o);

  input a;
  input b;
  input s;
  output o;
  assign o=(s==0)?b:a;

endmodule

module barrelLeft(i,s,o);      

	input[24:0] i;//25-bit Input line 
	input[4:0] s; //5 bit Shift magnitude
	output[24:0] o; //8-bit Output line 

	wire s1_1, s1_2, s1_3, s1_4, s1_5, s1_6, s1_7, s1_8, s1_9, s1_10, s1_11, s1_12, s1_13, s1_14, s1_15, s1_16, s1_17, s1_18, s1_19, s1_20, s1_21, s1_22, s1_23, s1_24, s1_25;
	wire s2_1, s2_2, s2_3, s2_4, s2_5, s2_6, s2_7, s2_8, s2_9, s2_10, s2_11, s2_12, s2_13, s2_14, s2_15, s2_16, s2_17, s2_18, s2_19, s2_20, s2_21, s2_22, s2_23, s2_24, s2_25;
	wire s3_1, s3_2, s3_3, s3_4, s3_5, s3_6, s3_7, s3_8, s3_9, s3_10, s3_11, s3_12, s3_13, s3_14, s3_15, s3_16, s3_17, s3_18, s3_19, s3_20, s3_21, s3_22, s3_23, s3_24, s3_25;
	wire s4_1, s4_2, s4_3, s4_4, s4_5, s4_6, s4_7, s4_8, s4_9, s4_10, s4_11, s4_12, s4_13, s4_14, s4_15, s4_16, s4_17, s4_18, s4_19, s4_20, s4_21, s4_22, s4_23, s4_24, s4_25;

	//stage 1
	mux m1(1'b0, i[0], s[0], s1_1);
	mux m2(i[0], i[1], s[0], s1_2);
	mux m3(i[1], i[2], s[0], s1_3);
	mux m4(i[2], i[3], s[0], s1_4);
	mux m5(i[3], i[4], s[0], s1_5);
	mux m6(i[4], i[5], s[0], s1_6);
	mux m7(i[5], i[6], s[0], s1_7);
	mux m8(i[6], i[7], s[0], s1_8);
	mux m9(i[7], i[8], s[0], s1_9);
	mux m10(i[8], i[9], s[0], s1_10);
	mux m11(i[9], i[10], s[0], s1_11);
	mux m12(i[10], i[11], s[0], s1_12);
	mux m13(i[11], i[12], s[0], s1_13);
	mux m14(i[12], i[13], s[0], s1_14);
	mux m15(i[13], i[14], s[0], s1_15);
	mux m16(i[14], i[15], s[0], s1_16);
	mux m17(i[15], i[16], s[0], s1_17);
	mux m18(i[16], i[17], s[0], s1_18);
	mux m19(i[17], i[18], s[0], s1_19);
	mux m20(i[18], i[19], s[0], s1_20);
	mux m21(i[19], i[20], s[0], s1_21);
	mux m22(i[20], i[21], s[0], s1_22);
	mux m23(i[21], i[22], s[0], s1_23);
	mux m24(i[22], i[23], s[0], s1_24);
	mux m24x(i[23], i[24], s[0], s1_25);

	//stage 2
	mux m25(1'b0, s1_1, s[1], s2_1);
	mux m26(1'b0, s1_2, s[1], s2_2);
	mux m27(s1_1, s1_3, s[1], s2_3);
	mux m28(s1_2, s1_4, s[1], s2_4);
	mux m29(s1_3, s1_5, s[1], s2_5);
	mux m30(s1_4, s1_6, s[1], s2_6);
	mux m31(s1_5, s1_7, s[1], s2_7);
	mux m32(s1_6, s1_8, s[1], s2_8);
	mux m33(s1_7, s1_9, s[1], s2_9);
	mux m34(s1_8, s1_10, s[1], s2_10);
	mux m35(s1_9, s1_11, s[1], s2_11);
	mux m36(s1_10, s1_12, s[1], s2_12);
	mux m37(s1_11, s1_13, s[1], s2_13);
	mux m38(s1_12, s1_14, s[1], s2_14);
	mux m39(s1_13, s1_15, s[1], s2_15);
	mux m40(s1_14, s1_16, s[1], s2_16);
	mux m41(s1_15, s1_17, s[1], s2_17);
	mux m42(s1_16, s1_18, s[1], s2_18);
	mux m43(s1_17, s1_19, s[1], s2_19);
	mux m44(s1_18, s1_20, s[1], s2_20);
	mux m45(s1_19, s1_21, s[1], s2_21);
	mux m46(s1_20, s1_22, s[1], s2_22);
	mux m47(s1_21, s1_23, s[1], s2_23);
	mux m48(s1_22, s1_24, s[1], s2_24);
	mux m48x(s1_23, s1_25, s[1], s2_25);

	//stage 3
	mux m49(1'b0, s2_1, s[2], s3_1);
	mux m50(1'b0, s2_2, s[2], s3_2);
	mux m51(1'b0, s2_3, s[2], s3_3);
	mux m52(1'b0, s2_4, s[2], s3_4);
	mux m53(s2_1, s2_5, s[2], s3_5);
	mux m54(s2_2, s2_6, s[2], s3_6);
	mux m55(s2_3, s2_7, s[2], s3_7);
	mux m56(s2_4, s2_8, s[2], s3_8);
	mux m57(s2_5, s2_9, s[2], s3_9);
	mux m58(s2_6, s2_10, s[2], s3_10);
	mux m59(s2_7, s2_11, s[2], s3_11);
	mux m60(s2_8, s2_12, s[2], s3_12);
	mux m61(s2_9, s2_13, s[2], s3_13);
	mux m62(s2_10, s2_14, s[2], s3_14);
	mux m63(s2_11, s2_15, s[2], s3_15);
	mux m64(s2_12, s2_16, s[2], s3_16);
	mux m65(s2_13, s2_17, s[2], s3_17);
	mux m66(s2_14, s2_18, s[2], s3_18);
	mux m67(s2_15, s2_19, s[2], s3_19);
	mux m68(s2_16, s2_20, s[2], s3_20);
	mux m69(s2_17, s2_21, s[2], s3_21);
	mux m70(s2_18, s2_22, s[2], s3_22);
	mux m71(s2_19, s2_23, s[2], s3_23);
	mux m72(s2_20, s2_24, s[2], s3_24);
	mux m72x(s2_21, s2_25, s[2], s3_25);

	//stage 4
	mux m73(1'b0, s3_1, s[3], s4_1);
	mux m74(1'b0, s3_2, s[3], s4_2);
	mux m75(1'b0, s3_3, s[3], s4_3);
	mux m76(1'b0, s3_4, s[3], s4_4);
	mux m77(1'b0, s3_5, s[3], s4_5);
	mux m78(1'b0, s3_6, s[3], s4_6);
	mux m79(1'b0, s3_7, s[3], s4_7);
	mux m80(1'b0, s3_8, s[3], s4_8);
	mux m81(s3_1, s3_9, s[3], s4_9);
	mux m82(s3_2, s3_10, s[3], s4_10);
	mux m83(s3_3, s3_11, s[3], s4_11);
	mux m84(s3_4, s3_12, s[3], s4_12);
	mux m85(s3_5, s3_13, s[3], s4_13);
	mux m86(s3_6, s3_14, s[3], s4_14);
	mux m87(s3_7, s3_15, s[3], s4_15);
	mux m88(s3_8, s3_16, s[3], s4_16);
	mux m89(s3_9, s3_17, s[3], s4_17);
	mux m90(s3_10, s3_18, s[3], s4_18);
	mux m91(s3_11, s3_19, s[3], s4_19);
	mux m92(s3_12, s3_20, s[3], s4_20);
	mux m93(s3_13, s3_21, s[3], s4_21);
	mux m94(s3_14, s3_22, s[3], s4_22);
	mux m95(s3_15, s3_23, s[3], s4_23);
	mux m96(s3_16, s3_24, s[3], s4_24);
	mux m96x(s3_17, s3_25, s[3], s4_25);

	//stage 5
	mux m97(1'b0, s4_1, s[4], o[0]);
	mux m98(1'b0, s4_2, s[4], o[1]);
	mux m99(1'b0, s4_3, s[4], o[2]);
	mux m100(1'b0, s4_4, s[4], o[3]);
	mux m101(1'b0, s4_5, s[4], o[4]);
	mux m102(1'b0, s4_6, s[4], o[5]);
	mux m103(1'b0, s4_7, s[4], o[6]);
	mux m104(1'b0, s4_8, s[4], o[7]);
	mux m105(1'b0, s4_9, s[4], o[8]);
	mux m106(1'b0, s4_10, s[4], o[9]);
	mux m107(1'b0, s4_11, s[4], o[10]);
	mux m108(1'b0, s4_12, s[4], o[11]);
	mux m109(1'b0, s4_13, s[4], o[12]);
	mux m110(1'b0, s4_14, s[4], o[13]);
	mux m111(1'b0, s4_15, s[4], o[14]);
	mux m112(1'b0, s4_16, s[4], o[15]);
	mux m113(s4_1, s4_17, s[4], o[16]);
	mux m114(s4_2, s4_18, s[4], o[17]);
	mux m115(s4_3, s4_19, s[4], o[18]);
	mux m116(s4_4, s4_20, s[4], o[19]);
	mux m117(s4_5, s4_21, s[4], o[20]);
	mux m118(s4_6, s4_22, s[4], o[21]);
	mux m119(s4_7, s4_23, s[4], o[22]);
	mux m120(s4_8, s4_24, s[4], o[23]);
	mux m120x(s4_9, s4_25, s[4], o[24]);

endmodule

module barrelRight(i,s,o);   

	input[23:0] i;//24-bit Input line 
	input[4:0] s; //5 bit Shift magnitude
	output[23:0] o; //8-bit Output line 

	wire s1_1, s1_2, s1_3, s1_4, s1_5, s1_6, s1_7, s1_8, s1_9, s1_10, s1_11, s1_12, s1_13, s1_14, s1_15, s1_16, s1_17, s1_18, s1_19, s1_20, s1_21, s1_22, s1_23, s1_24;
	wire s2_1, s2_2, s2_3, s2_4, s2_5, s2_6, s2_7, s2_8, s2_9, s2_10, s2_11, s2_12, s2_13, s2_14, s2_15, s2_16, s2_17, s2_18, s2_19, s2_20, s2_21, s2_22, s2_23, s2_24;
	wire s3_1, s3_2, s3_3, s3_4, s3_5, s3_6, s3_7, s3_8, s3_9, s3_10, s3_11, s3_12, s3_13, s3_14, s3_15, s3_16, s3_17, s3_18, s3_19, s3_20, s3_21, s3_22, s3_23, s3_24;
	wire s4_1, s4_2, s4_3, s4_4, s4_5, s4_6, s4_7, s4_8, s4_9, s4_10, s4_11, s4_12, s4_13, s4_14, s4_15, s4_16, s4_17, s4_18, s4_19, s4_20, s4_21, s4_22, s4_23, s4_24;

	//stage 1
	mux m1(i[1], i[0], s[0], s1_1);
	mux m2(i[2], i[1], s[0], s1_2);
	mux m3(i[3], i[2], s[0], s1_3);
	mux m4(i[4], i[3], s[0], s1_4);
	mux m5(i[5], i[4], s[0], s1_5);
	mux m6(i[6], i[5], s[0], s1_6);
	mux m7(i[7], i[6], s[0], s1_7);
	mux m8(i[8], i[7], s[0], s1_8);
	mux m9(i[9], i[8], s[0], s1_9);
	mux m10(i[10], i[9], s[0], s1_10);
	mux m11(i[11], i[10], s[0], s1_11);
	mux m12(i[12], i[11], s[0], s1_12);
	mux m13(i[13], i[12], s[0], s1_13);
	mux m14(i[14], i[13], s[0], s1_14);
	mux m15(i[15], i[14], s[0], s1_15);
	mux m16(i[16], i[15], s[0], s1_16);
	mux m17(i[17], i[16], s[0], s1_17);
	mux m18(i[18], i[17], s[0], s1_18);
	mux m19(i[19], i[18], s[0], s1_19);
	mux m20(i[20], i[19], s[0], s1_20);
	mux m21(i[21], i[20], s[0], s1_21);
	mux m22(i[22], i[21], s[0], s1_22);
	mux m23(i[23], i[22], s[0], s1_23);
	mux m24(1'b0, i[23], s[0], s1_24);

	//stage 2
	mux m25(s1_3, s1_1, s[1], s2_1);
	mux m26(s1_4, s1_2, s[1], s2_2);
	mux m27(s1_5, s1_3, s[1], s2_3);
	mux m28(s1_6, s1_4, s[1], s2_4);
	mux m29(s1_7, s1_5, s[1], s2_5);
	mux m30(s1_8, s1_6, s[1], s2_6);
	mux m31(s1_9, s1_7, s[1], s2_7);
	mux m32(s1_10, s1_8, s[1], s2_8);
	mux m33(s1_11, s1_9, s[1], s2_9);
	mux m34(s1_12, s1_10, s[1], s2_10);
	mux m35(s1_13, s1_11, s[1], s2_11);
	mux m36(s1_14, s1_12, s[1], s2_12);
	mux m37(s1_15, s1_13, s[1], s2_13);
	mux m38(s1_16, s1_14, s[1], s2_14);
	mux m39(s1_17, s1_15, s[1], s2_15);
	mux m40(s1_18, s1_16, s[1], s2_16);
	mux m41(s1_19, s1_17, s[1], s2_17);
	mux m42(s1_20, s1_18, s[1], s2_18);
	mux m43(s1_21, s1_19, s[1], s2_19);
	mux m44(s1_22, s1_20, s[1], s2_20);
	mux m45(s1_23, s1_21, s[1], s2_21);
	mux m46(s1_24, s1_22, s[1], s2_22);
	mux m47(1'b0, s1_23, s[1], s2_23);
	mux m48(1'b0, s1_24, s[1], s2_24);

	//stage 3
	mux m49(s2_5, s2_1, s[2], s3_1);
	mux m50(s2_6, s2_2, s[2], s3_2);
	mux m51(s2_7, s2_3, s[2], s3_3);
	mux m52(s2_8, s2_4, s[2], s3_4);
	mux m53(s2_9, s2_5, s[2], s3_5);
	mux m54(s2_10, s2_6, s[2], s3_6);
	mux m55(s2_11, s2_7, s[2], s3_7);
	mux m56(s2_12, s2_8, s[2], s3_8);
	mux m57(s2_13, s2_9, s[2], s3_9);
	mux m58(s2_14, s2_10, s[2], s3_10);
	mux m59(s2_15, s2_11, s[2], s3_11);
	mux m60(s2_16, s2_12, s[2], s3_12);
	mux m61(s2_17, s2_13, s[2], s3_13);
	mux m62(s2_18, s2_14, s[2], s3_14);
	mux m63(s2_19, s2_15, s[2], s3_15);
	mux m64(s2_20, s2_16, s[2], s3_16);
	mux m65(s2_21, s2_17, s[2], s3_17);
	mux m66(s2_22, s2_18, s[2], s3_18);
	mux m67(s2_23, s2_19, s[2], s3_19);
	mux m68(s2_24, s2_20, s[2], s3_20);
	mux m69(1'b0, s2_21, s[2], s3_21);
	mux m70(1'b0, s2_22, s[2], s3_22);
	mux m71(1'b0, s2_23, s[2], s3_23);
	mux m72(1'b0, s2_24, s[2], s3_24);

	//stage 4
	mux m73(s3_9, s3_1, s[3], s4_1);
	mux m74(s3_10, s3_2, s[3], s4_2);
	mux m75(s3_11, s3_3, s[3], s4_3);
	mux m76(s3_12, s3_4, s[3], s4_4);
	mux m77(s3_13, s3_5, s[3], s4_5);
	mux m78(s3_14, s3_6, s[3], s4_6);
	mux m79(s3_15, s3_7, s[3], s4_7);
	mux m80(s3_16, s3_8, s[3], s4_8);
	mux m81(s3_17, s3_9, s[3], s4_9);
	mux m82(s3_18, s3_10, s[3], s4_10);
	mux m83(s3_19, s3_11, s[3], s4_11);
	mux m84(s3_20, s3_12, s[3], s4_12);
	mux m85(s3_21, s3_13, s[3], s4_13);
	mux m86(s3_22, s3_14, s[3], s4_14);
	mux m87(s3_23, s3_15, s[3], s4_15);
	mux m88(s3_24, s3_16, s[3], s4_16);
	mux m89(1'b0, s3_17, s[3], s4_17);
	mux m90(1'b0, s3_18, s[3], s4_18);
	mux m91(1'b0, s3_19, s[3], s4_19);
	mux m92(1'b0, s3_20, s[3], s4_20);
	mux m93(1'b0, s3_21, s[3], s4_21);
	mux m94(1'b0, s3_22, s[3], s4_22);
	mux m95(1'b0, s3_23, s[3], s4_23);
	mux m96(1'b0, s3_24, s[3], s4_24);

	//stage 5
	mux m97(s4_17, s4_1, s[4], o[0]);
	mux m98(s4_18, s4_2, s[4], o[1]);
	mux m99(s4_19, s4_3, s[4], o[2]);
	mux m100(s4_20, s4_4, s[4], o[3]);
	mux m101(s4_21, s4_5, s[4], o[4]);
	mux m102(s4_22, s4_6, s[4], o[5]);
	mux m103(s4_23, s4_7, s[4], o[6]);
	mux m104(s4_24, s4_8, s[4], o[7]);
	mux m105(1'b0, s4_9, s[4], o[8]);
	mux m106(1'b0, s4_10, s[4], o[9]);
	mux m107(1'b0, s4_11, s[4], o[10]);
	mux m108(1'b0, s4_12, s[4], o[11]);
	mux m109(1'b0, s4_13, s[4], o[12]);
	mux m110(1'b0, s4_14, s[4], o[13]);
	mux m111(1'b0, s4_15, s[4], o[14]);
	mux m112(1'b0, s4_16, s[4], o[15]);
	mux m113(1'b0, s4_17, s[4], o[16]);
	mux m114(1'b0, s4_18, s[4], o[17]);
	mux m115(1'b0, s4_19, s[4], o[18]);
	mux m116(1'b0, s4_20, s[4], o[19]);
	mux m117(1'b0, s4_21, s[4], o[20]);
	mux m118(1'b0, s4_22, s[4], o[21]);
	mux m119(1'b0, s4_23, s[4], o[22]);
	mux m120(1'b0, s4_24, s[4], o[23]);

endmodule